module class(
		input a,
		output b
		)

assign b = a;

endmodule